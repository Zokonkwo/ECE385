module alu (input logic [15:0] sr2mux, sr1out, 
            input logic [2:0] aluk,
            output logic [15:0] alu_out);



  
endmodule
