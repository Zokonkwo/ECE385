module bit3__mux_2_1()
