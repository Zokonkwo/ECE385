module reg_file2()
endmodule
