module decoder (input logic [15:0] ir_in,
                input logic clk,
                output logic [15:0] decoder_out);

endmodule
