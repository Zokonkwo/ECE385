module nzp (input logic ld_cc
           );

endmodule 
