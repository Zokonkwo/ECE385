module decoder (input logic [15:0] ir_in,
                output logic [15:0] decoder_out);

endmodule
